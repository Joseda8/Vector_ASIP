module plus_1 (input logic  [31:0] a, output logic [31:0] s);
	  
	assign s = a + 1;
	
endmodule 