module datapath(clk, rst, instr_in, wr_pixels, algorithm, wr_wom, vec_func, pc, instr_out);

	input logic clk, rst, wr_pixels, algorithm, wr_wom, vec_func;
	input logic [29:0] instr_in;
	
	output logic [29:0] instr_out;
	output logic [31:0] pc;
	
	
	
	


endmodule
